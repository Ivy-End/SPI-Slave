`ifndef __UTILS__
`define __UTILS__

class Utils;
    extern task WaveformDump(string waveformName);
endclass

task Utils::WaveformDump(string waveformName);
endtask

`endif